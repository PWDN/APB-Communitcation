module apb_slave_exe_w47(i_PDATA,
                        i_PRESETn,
                        i_PADDR,
                        i_PSEL,
                        i_PENABLE,
                        i_PWDATA,
                        o_READY,
                        o_PRDATA,
                        o_PSLVERR);



endmodule
