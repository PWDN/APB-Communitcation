`ifndef PARAMS_DEFINE
`define PARAMS_DEFINE

`define DATA_WIDTH 4
`define ADDR_WIDTH 16
`define SEL_WIDTH 16

`define CLK_STEP 3
`endif
