`ifndef PARAMS_DEFINE
`define PARAMS_DEFINE

`define DATA_WIDTH 8
`define ADDR_WIDTH 16
`define SEL_WIDTH 2

`define CLK_STEP 3

`define ARG_WIDTH 3
`define STATUS_WIDTH 4

`endif
